<?xml version="1.0" encoding="UTF-8"?>
<svg version="1.1" xmlns="http://www.w3.org/2000/svg" width="512" height="512" viewBox="25 30 465 465">
<path d="M0 0 C1.32268101 -0.00551503 1.32268101 -0.00551503 2.67208284 -0.01114148 C5.63282978 -0.02217228 8.59354162 -0.02602117 11.55430603 -0.02983093 C13.67495332 -0.03609611 15.79559952 -0.04274296 17.91624451 -0.04974365 C24.88665503 -0.07078256 31.85706576 -0.0811469 38.82749939 -0.09111023 C41.22817433 -0.09515806 43.62884915 -0.09927499 46.02952385 -0.10346031 C57.30999606 -0.12251277 68.59046173 -0.13674286 79.87094694 -0.14507228 C92.88516032 -0.15484082 105.89920344 -0.18115027 118.91335684 -0.22157317 C128.9763726 -0.25175501 139.03933963 -0.26654319 149.10239977 -0.26985329 C155.11052945 -0.27220169 161.11847725 -0.28113492 167.1265583 -0.30631447 C172.78270033 -0.32963573 178.43854125 -0.33381195 184.09471893 -0.32355309 C186.16547333 -0.32305858 188.23624275 -0.32935369 190.30695152 -0.34310913 C205.91491661 -0.44095049 218.75418748 0.93942476 230.55015564 12.25263977 C240.50228887 22.92088591 242.65654248 33.42538786 242.64537048 47.70674133 C242.65208771 48.94684464 242.65880493 50.18694794 242.66572571 51.46463013 C242.68140887 54.8471611 242.68807725 58.22944642 242.68935728 61.61199665 C242.6907848 63.73147683 242.69506575 65.85093172 242.70035172 67.97040558 C242.71882312 75.3823712 242.72702611 82.79426518 242.72544861 90.20625305 C242.72424853 97.08637944 242.74533182 103.96619146 242.77693594 110.84623837 C242.80319616 116.77691391 242.81381182 122.7074874 242.81253779 128.63822055 C242.81203094 132.16981255 242.81755891 135.70112494 242.83889389 139.23265839 C242.86208407 143.17856817 242.85269603 147.12405605 242.84068298 151.07002258 C242.851922 152.22055618 242.86316101 153.37108978 242.8747406 154.55648804 C242.76853929 168.36004418 238.1151777 179.50244665 228.25718689 189.21357727 C219.24495294 196.78647077 211.09497234 199.14717102 199.35484314 199.14717102 C199.35484314 217.95717102 199.35484314 236.76717102 199.35484314 256.14717102 C191.53813207 249.44713296 191.53813207 249.44713296 188.21604919 244.92973328 C164.04219654 212.94804075 164.04219654 212.94804075 128.88340759 196.59978104 C109.96876608 194.03938814 90.6048192 195.15253235 71.62084198 196.32661986 C62.02806507 196.91055922 52.42988534 197.16283407 42.82359314 197.41279602 C39.43065864 197.50256356 36.03779732 197.59453174 32.64500427 197.6894989 C31.41256131 197.72392233 31.41256131 197.72392233 30.15522051 197.75904119 C24.55890612 197.92440956 18.97104297 198.17720955 13.38011169 198.47032166 C11.16821415 198.57837967 8.95625225 198.68501916 6.74427032 198.79133415 C4.72519542 198.89571295 2.70739145 199.02384548 0.68974304 199.15289307 C-10.91994375 199.70791362 -19.6191287 196.4461974 -28.64515686 189.14717102 C-36.06331116 182.29140387 -42.2243206 173.0086767 -42.77937794 162.63983059 C-42.78365142 161.69176572 -42.7879249 160.74370085 -42.79232788 159.76690674 C-42.79948318 158.67505066 -42.80663849 157.58319458 -42.81401062 156.45825195 C-42.81804398 154.66832573 -42.81804398 154.66832573 -42.82215881 152.84223938 C-42.82873001 151.58160675 -42.83530121 150.32097412 -42.84207153 149.0221405 C-42.86307233 144.84377811 -42.87347334 140.66541554 -42.88343811 136.48701477 C-42.8874878 135.04472396 -42.89160478 133.60243333 -42.89578819 132.1601429 C-42.91483476 125.37968452 -42.92906432 118.59923697 -42.93740016 111.818757 C-42.94715705 104.01269886 -42.97343801 96.20692545 -43.01390105 88.40096754 C-43.04415671 82.35490278 -43.05887813 76.30891918 -43.06218117 70.26278025 C-43.0645218 66.65792696 -43.07335155 63.05337801 -43.09864235 59.44860649 C-43.12646239 55.41817998 -43.12206326 51.38838109 -43.11512756 47.35786438 C-43.12793762 46.17874985 -43.14074768 44.99963531 -43.15394592 43.78479004 C-43.0741148 31.00509576 -38.65604438 20.48069938 -30.14515686 11.02217102 C-21.81451433 2.96179743 -11.2428988 -0.0025119 0 0 Z " fill="#000000" transform="translate(241.64515686035156,184.8528289794922)"/>
<path d="M0 0 C0.85743488 -0.00297112 1.71486977 -0.00594224 2.59828752 -0.0090034 C5.4706812 -0.01767304 8.34303312 -0.0191972 11.21543884 -0.02069092 C13.27549834 -0.02532041 15.33555698 -0.03034525 17.39561462 -0.03573608 C22.99305287 -0.0488516 28.59047913 -0.05530368 34.18793035 -0.05974674 C37.68749798 -0.06267954 41.18706235 -0.06678479 44.68662834 -0.07125092 C55.64300206 -0.08492516 66.5993683 -0.09459152 77.55574995 -0.09845281 C90.18957023 -0.10293002 102.82328213 -0.12046268 115.45706946 -0.1494534 C125.23052759 -0.17109928 135.00395531 -0.18115868 144.77743715 -0.18249393 C150.61060945 -0.1835401 156.44367986 -0.18940767 162.27682686 -0.20731354 C167.76879556 -0.22384386 173.26058633 -0.22592563 178.75257111 -0.21717453 C180.76162379 -0.21640674 182.77068624 -0.22071255 184.77971458 -0.23063278 C201.23647894 -0.30708776 214.97482152 0.64902876 227.75816345 12.21075439 C236.2066098 21.0389062 239.64319394 30.83949493 239.5667572 42.84356689 C239.56463478 44.10025177 239.56463478 44.10025177 239.56246948 45.38232422 C239.55688293 48.05173347 239.54433289 50.7210581 239.53160095 53.39044189 C239.52658421 55.20294068 239.52202161 57.01544079 239.51792908 58.82794189 C239.50691789 63.26547438 239.4896625 67.7029438 239.46910095 72.14044189 C238.5104715 72.14630814 237.55184204 72.15217438 236.56416321 72.15821838 C227.47378832 72.21574746 218.38364575 72.28866286 209.29350853 72.37615681 C204.62158856 72.42064338 199.94975146 72.45994561 195.2776947 72.48687744 C190.75820854 72.51312926 186.23904506 72.5536812 181.71976089 72.60362816 C180.00648171 72.62015047 178.29314691 72.63175488 176.57979965 72.6380558 C154.13944784 72.72882853 134.67954565 77.85594269 117.71910095 93.32794189 C102.39193991 109.87517546 98.24747671 130.16768505 98.05503845 152.09356689 C98.03627528 153.48890257 98.01669829 154.88422751 97.99635315 156.27954102 C97.94556846 159.90923663 97.90566 163.53896883 97.86820984 167.16882324 C97.8278287 170.88991946 97.77689415 174.61087067 97.72691345 178.33184814 C97.63079189 185.60127902 97.54618857 192.87078157 97.46910095 200.14044189 C96.45976501 199.87747314 95.45042908 199.61450439 94.4105072 199.34356689 C81.20347643 196.27543126 67.00229435 195.2460015 54.46910095 201.14044189 C33.54932225 214.46514226 16.56240484 236.47433363 0.42597961 255.02119446 C-0.54267532 256.07022194 -0.54267532 256.07022194 -1.53089905 257.14044189 C-1.86089905 257.14044189 -2.19089905 257.14044189 -2.53089905 257.14044189 C-2.53089905 238.33044189 -2.53089905 219.52044189 -2.53089905 200.14044189 C-6.16089905 199.81044189 -9.79089905 199.48044189 -13.53089905 199.14044189 C-25.89688265 195.11777253 -35.24796928 187.76096882 -41.34339905 176.14044189 C-45.45364176 167.83578769 -45.82546263 159.93690901 -45.80555725 150.84039307 C-45.81066818 149.62794418 -45.81577911 148.4154953 -45.82104492 147.16630554 C-45.83251711 143.86027782 -45.83502182 140.55450184 -45.83248162 137.24847198 C-45.83140655 134.4779572 -45.83630906 131.70746515 -45.84108704 128.93695527 C-45.8521572 122.39400815 -45.85263412 115.85111845 -45.84657288 109.3081665 C-45.84053871 102.58371194 -45.85283554 95.85946692 -45.87414294 89.13504809 C-45.89182441 83.33942028 -45.89774993 77.54385876 -45.8945052 71.74820501 C-45.89270213 68.29662421 -45.89522969 64.8451928 -45.90921974 61.3936367 C-45.92426239 57.53856738 -45.91477099 53.68375971 -45.9032135 49.82867432 C-45.91085724 48.70259766 -45.91850098 47.576521 -45.92637634 46.4163208 C-45.83788841 32.9968369 -42.06598183 20.8922311 -32.53089905 11.14044189 C-22.69668333 3.33954314 -12.44326673 -0.01350705 0 0 Z " fill="#000000" transform="translate(73.53089904785156,84.85955810546875)"/>
</svg>
